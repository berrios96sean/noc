// parameters.sv
`ifndef PARAMETERS_SV
`define PARAMETERS_SV

// Define your parameters here
parameter int ROWS = 2;
parameter int COLUMNS = 2;

`endif // PARAMETERS_SV
